
module controller(
    input clk, reset,

    // Decode stage control signals
    input [6:0] opD,
    input [2:0] funct3D,
    input funct7b5D,
    output [2:0] ImmSrcD,

    // Execute stage control signals
    input FlushE,
    input [3:0] FlagE,
    output PCSrcE, // for datapath and Hazard Unit
    output [3:0] ALUControlE,
    output ALUSrcAE,
    output ALUSrcBE, // for lui
    output [1:0] PCSrcSelE, // for jalr
    output ResultSrcEb0, // for Hazard Unit

    // Memory stage control signals
    output MemWriteM,
    output RegWriteM, // for Hazard Unit

    // Writeback stage control signals
    output RegWriteW, // for datapath and Hazard Unit
    output [1:0] ResultSrcW,
    
    output [2:0]LoadType,
    output [1:0]StoreType
);

    // pipelined control signals
    wire RegWriteD, RegWriteE;
    wire [1:0] ResultSrcD, ResultSrcE, ResultSrcM;
    wire MemWriteD, MemWriteE;
    wire JumpD, JumpE;
    wire BranchD, BranchE;
    wire [1:0] ALUOpD;
    wire [3:0] ALUControlD;
    wire ALUSrcAD;
    wire ALUSrcBD; // for lui
    wire takenE;
    wire [2:0] funct3E;
    wire JALRD, JALRE; // for jalr
    wire [2:0] LoadTypeD, LoadTypeE, LoadTypeM;
    wire [1:0] StoreTypeD, StoreTypeE, StoreTypeM;
    // Decode stage logic
    maindec md(
        .op(opD),
        .ResultSrc(ResultSrcD),
        .MemWrite(MemWriteD),
        .Branch(BranchD),
        .ALUSrcA(ALUSrcAD),
        .ALUSrcB(ALUSrcBD),
        .RegWrite(RegWriteD),
        .Jump(JumpD),
        .JALR(JALRD),
        .ImmSrc(ImmSrcD),
        .ALUOp(ALUOpD)
    );
    aludec ad(
        .op5(opD[5]),
        .funct3(funct3D),
        .funct7b5(funct7b5D),
        .ALUOp(ALUOpD),
        .ALUControl(ALUControlD)
    );
  loadstoreunit lsu(.opcode(opD),.funct3(funct3D),.LoadType(LoadTypeD),.StoreType(StoreTypeD));
    
    // Execute stage pipeline control register and logic
   floprc #(21) controlregE( // +5 for 3+2 bits
    .clk(clk),
    .reset(reset),
    .clear(FlushE),
    .d({RegWriteD, ResultSrcD, MemWriteD, JumpD, BranchD, ALUControlD, ALUSrcAD, ALUSrcBD, funct3D, JALRD, LoadTypeD, StoreTypeD}),
    .q({RegWriteE, ResultSrcE, MemWriteE, JumpE, BranchE, ALUControlE, ALUSrcAE, ALUSrcBE, funct3E, JALRE, LoadTypeE, StoreTypeE})
);
    
    
    branchunit bu(
        .Branch (BranchE),   // From pipelined control register
        .Flags  (FlagE),     // From datapath/ALU
        .funct3 (funct3E),   // Pipelined from Decode stage
        .taken  (takenE)
    );

    assign PCSrcE = takenE | JumpE;
    assign PCSrcSelE = JALRE        ? 2'b10 :
                   (takenE | JumpE) ? 2'b01 :
                   2'b00;
    assign ResultSrcEb0 = ResultSrcE[0];

    // Memory stage pipeline control register
    flopr #(9) controlregM(.clk(clk),
    .reset(reset),
    .d({RegWriteE, ResultSrcE, MemWriteE, LoadTypeE, StoreTypeE}),
    .q({RegWriteM, ResultSrcM, MemWriteM, LoadTypeM, StoreTypeM}));
     assign LoadType  = LoadTypeM;
     assign StoreType = StoreTypeM;

    // Writeback stage pipeline control register
    flopr #(3) controlregW(
        .clk(clk),
        .reset(reset),
        .d({RegWriteM, ResultSrcM}),
        .q({RegWriteW, ResultSrcW})
    );

endmodule